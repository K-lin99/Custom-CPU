library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity icache is
port(   	i_cache_address	 : in  std_logic_vector(4 downto 0);
		data_out         : out std_logic_vector(31 downto 0)		);
end icache ;

architecture rtl of icache is
begin

	with i_cache_address select                      --  rd|rt,rs rt
	data_out <= "00100000000000110000000000000000" when "00000",  
				"00100000000000010000000000000000" when "00001", 
				"00100000000000100000000000000101" when "00010", 
				"00000000001000100000100000100000" when "00011", 
				"00100000010000101111111111111111" when "00100", 
				"00010000010000110000000000000001" when "00101", 
				"00001000000000000000000000000011" when "00110", 
				"10101100000000010000000000000000" when "00111", 
				"10001100000001000000000000000000" when "01000", 
				"00110000100001000000000000001010" when "01001", 
				"00110100100001000000000000000001" when "01010", 
				"00111000100001000000000000001011" when "01011", 
				"00111000100001000000000000000000" when "01100", 
				"00000000000000000000000000000000" when others; 
end;

